** Profile: "SCHEMATIC1-ac-sweep"  [ C:\Users\Usuario_UMA\Downloads\CREATIVA\CREATIVA\CREATIVA\MESA_DE_MEZCLAS-PSpiceFiles\SCHEMATIC1\ac-sweep.sim ] 

** Creating circuit file "ac-sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Usuario_UMA\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC OCT 100 20 20000
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
